----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/20/2024 02:42:50 PM
-- Design Name: 
-- Module Name: complex_comp - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity complex_comp is
    generic ( nbits : integer := 4);
    Port ( a : in STD_LOGIC_vector(nbits-1 downto 0);
           b : in std_logic_vector(nbits-1 downto 0);
           o : out STD_LOGIC);
end complex_comp;

architecture Behavioral of complex_comp is

begin
process(a,b)
    begin
    if(unsigned(a) < unsigned(b)) then
        o <= '1';
        else
        o <= '0';
        end if;
end process;

end Behavioral;
